
module TEST_OY_CPU (
	clk_clk);	

	input		clk_clk;
endmodule
